module FIFOBuffer (q
    
);
    
endmodule