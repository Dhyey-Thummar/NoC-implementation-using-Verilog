module FIFOBuffer (q,k
    
);
    
endmodule