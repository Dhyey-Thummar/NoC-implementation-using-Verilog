module FIFOBuffer (
    
);
    
endmodule